CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files (x86)\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9961490 0
0
6 Title:
5 Name:
0
0
0
10
9 Resistor~
219 768 274 0 3 5
0 2 3 -1
0
0 0 864 90
4 1.1M
21 4 49 12
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3472 0 0
2
41716.7 0
0
10 Polar Cap~
219 732 271 0 2 5
0 3 2
0
0 0 832 270
5 2.2uF
-44 10 -9 18
2 C2
14 -6 28 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9998 0 0
2
41716.7 0
0
7 Op Amp~
219 638 240 0 1 7
0 0
0
0 0 832 0
5 IDEAL
-18 -25 17 -17
2 U2
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 0 0 0 0
1 U
3536 0 0
2
41716.7 0
0
7 Ground~
168 439 116 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
41716.7 0
0
9 Resistor~
219 480 202 0 2 5
0 5 6
0
0 0 864 180
3 22K
-11 -14 10 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3835 0 0
2
41716.7 0
0
9 Resistor~
219 439 168 0 2 5
0 5 6
0
0 0 864 90
3 100
7 0 28 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3670 0 0
2
41716.7 0
0
7 Op Amp~
219 476 246 0 1 7
0 0
0
0 0 832 0
5 IDEAL
-18 -25 17 -17
2 U1
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 0 0 0 0
1 U
5616 0 0
2
41716.7 0
0
7 Ground~
168 746 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9323 0 0
2
5.89653e-315 0
0
6 Diode~
219 680 240 0 2 5
0 4 3
0
0 0 832 0
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
317 0 0
2
5.89653e-315 0
0
9 Resistor~
219 566 246 0 2 5
0 5 6
0
0 0 864 0
3 100
-9 -11 12 -3
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3108 0 0
2
5.89653e-315 0
0
14
1 0 0 0 0 0 0 8 0 0 2 2
746 309
746 300
2 1 0 0 0 0 0 2 1 0 0 4
731 278
731 300
768 300
768 292
2 0 0 0 0 0 0 1 0 0 6 2
768 256
768 240
1 0 0 0 0 0 0 2 0 0 6 2
731 261
731 240
2 0 0 0 0 0 0 3 0 0 6 5
620 234
608 234
608 180
707 180
707 240
2 0 0 0 0 0 0 9 0 0 0 2
690 240
787 240
1 3 0 0 0 0 0 5 7 0 0 4
498 202
517 202
517 246
494 246
2 1 0 0 0 0 0 6 4 0 0 2
439 150
439 124
2 0 0 0 0 0 0 5 0 0 10 2
462 202
439 202
2 1 0 0 0 0 0 7 6 0 0 3
458 240
439 240
439 186
0 1 0 0 0 0 0 0 7 0 0 2
363 252
458 252
0 1 0 0 0 0 0 0 10 7 0 3
517 245
517 246
548 246
3 1 4 0 0 4224 0 3 9 0 0 2
656 240
670 240
2 1 6 0 0 4224 0 10 3 0 0 2
584 246
620 246
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
777 221 820 245
782 225 814 241
4 Vout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
369 235 404 259
374 239 398 255
3 Vin
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
